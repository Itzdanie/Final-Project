module tb ();




endmodule